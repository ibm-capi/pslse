//
// Copyright 2014 International Business Machines
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

`timescale 1ns / 1ns

module top (
  output          breakpoint
);

   import "DPI-C" function void psl_bfm_init( );
   import "DPI-C" function void set_simulation_time(input [0:63] simulationTime);
   import "DPI-C" function void get_simuation_error(inout simulationError);
   import "DPI-C" function void psl_bfm( input ha_pclock, 
             inout           ha_jval_top, 
             inout  [0:7]    ha_jcom_top, 
             inout           ha_jcompar_top, 
             inout  [0:63]   ha_jea_top,
	     inout           ha_jeapar_top, 
             input           ah_jrunning_top,  
             input           ah_jdone_top,
	     input           ah_jcack_top, 
             input  [0:63]   ah_jerror_top, 
             input  [0:3]    ah_brlat_top,  
//             input           ah_jyield,
	     input           ah_tbreq_top, 
             input           ah_paren_top, 
             inout           ha_mmval_top,
             inout           ha_mmcfg_top, 
             inout           ha_mmrnw_top, 
             inout           ha_mmdw_top,
             inout  [0:23]   ha_mmad_top, 
             inout           ha_mmadpar_top, 
             inout  [0:63]   ha_mmdata_top, 
             inout           ha_mmdatapar_top,
             input           ah_mmack_top, 
             input [0:63]    ah_mmdata_top, 
             input           ah_mmdatapar_top,
             inout  [0:7]    ha_croom_top,
             input           ah_cvalid_top, 
             input  [0:7]    ah_ctag_top, 
             input           ah_ctagpar_top, 
             input  [0:12]   ah_com_top, 
             input           ah_compar_top, 
             input  [0:2]    ah_cabt_top, 
             input  [0:63]   ah_cea_top, 
             input           ah_ceapar_top, 
             input  [0:15]   ah_cch_top, 
             input  [0:11]   ah_csize_top, 
             input  [0:3]    ah_cpagesize_top, 
             inout           ha_brvalid_top, 
             inout  [0:7]    ha_brtag_top, 
             inout           ha_brtagpar_top, 
             input [0:1023]  ah_brdata_top, 
             input [0:15]    ah_brpar_top, 
             input           ah_brvalid_top, 
             input [0:7]     ah_brtag_top,
             inout           ha_bwvalid_top, 
             inout  [0:7]    ha_bwtag_top, 		// 8 bits
             inout           ha_bwtagpar_top,
             inout  [0:1023] ha_bwdata_top, 		// 1024 bits
             inout  [0:15]   ha_bwpar_top,	// 16 bits
             inout           ha_rvalid_top, 
             inout  [0:7]    ha_rtag_top, 		// 8 bits
             inout           ha_rtagpar_top,
             inout  [0:8]    ha_rditag_top,
             inout           ha_rditagpar_top,
             inout  [0:7]    ha_response_top, 		// 8 bits
             inout  [0:7]    ha_response_ext_top, 	// 8 bits
             inout  [0:3]    ha_rpagesize_top, 		// 4 bits
             inout  [0:1]    ha_rcachestate_top, 	// 2 bits
             inout  [0:12]   ha_rcachepos_top, 		// 13 bits
             inout  [0:8]    ha_rcredits_top,		// 9 bits
             input           d0h_dvalid_top,
             input  [0:9]    d0h_req_utag_top,
             input  [0:8]    d0h_req_itag_top,
             input  [0:2]    d0h_dtype_top,
             input  [0:9]    d0h_dsize_top,
             input  [0:1023] d0h_ddata_top,
             input  [0:5]    d0h_datomic_op_top,
             input           d0h_datomic_le_top,
	     inout           hd0_sent_utag_valid_top, 
	     inout  [0:9]    hd0_sent_utag_top, 
	     inout  [0:2]    hd0_sent_utag_sts_top, 
	     inout           hd0_cpl_valid_top, 
	     inout  [0:9]    hd0_cpl_utag_top, 
	     inout  [0:2]    hd0_cpl_type_top, 
	     inout  [0:9]    hd0_cpl_size_top, 
	     inout  [0:9]    hd0_cpl_laddr_top, 
	     inout  [0:9]    hd0_cpl_byte_count_top, 
             inout  [0:1023] hd0_cpl_data_top,
             input           d1h_dvalid_top,
             input  [0:9]    d1h_req_utag_top,
             input  [0:8]    d1h_req_itag_top,
             input  [0:2]    d1h_dtype_top,
             input  [0:9]    d1h_dsize_top,
             input  [0:1023] d1h_ddata_top,
             input  [0:5]    d1h_datomic_op_top,
             input           d1h_datomic_le_top,
	     inout           hd1_sent_utag_valid_top, 
	     inout  [0:9]    hd1_sent_utag_top, 
	     inout  [0:2]    hd1_sent_utag_sts_top, 
	     inout           hd1_cpl_valid_top, 
	     inout  [0:9]    hd1_cpl_utag_top, 
	     inout  [0:2]    hd1_cpl_type_top, 
	     inout  [0:9]    hd1_cpl_size_top, 
	     inout  [0:9]    hd1_cpl_laddr_top, 
	     inout  [0:9]    hd1_cpl_byte_count_top, 
             inout  [0:1023] hd1_cpl_data_top
             );
  // Input
  reg    [0:7]    ha_croom_top;
  reg             ha_brvalid_top;
  reg    [0:7]    ha_brtag_top;
  reg             ha_brtagpar_top;
  reg             ha_bwvalid_top;
  reg    [0:7]    ha_bwtag_top;
  reg             ha_bwtagpar_top;
  reg    [0:1023] ha_bwdata_top;
  reg    [0:15]   ha_bwpar_top;
  reg             ha_rvalid_top;
  reg    [0:7]    ha_rtag_top;
  reg             ha_rtagpar_top;
  reg    [0:8]    ha_rditag_top;
  reg             ha_rditagpar_top;
  reg    [0:7]    ha_response_top;
  reg    [0:7]    ha_response_ext_top;
  reg    [0:3]    ha_rpagesize_top;
  reg    [0:1]    ha_rcachestate_top;
  reg    [0:12]   ha_rcachepos_top;
  reg    [0:8]    ha_rcredits_top;
  reg             ha_mmval_top;
  reg             ha_mmcfg_top;
  reg             ha_mmrnw_top;
  reg             ha_mmdw_top;
  reg    [0:23]   ha_mmad_top;
  reg             ha_mmadpar_top;
  reg    [0:63]   ha_mmdata_top;
  reg             ha_mmdatapar_top;
  reg             ha_jval_top;
  reg    [0:7]    ha_jcom_top;
  reg             ha_jcompar_top;
  reg    [0:63]   ha_jea_top;
  reg             ha_jeapar_top;
  reg             ha_pclock;
  reg             hd0_sent_utag_valid_top;
  reg    [0:9]    hd0_sent_utag_top;
  reg    [0:2]    hd0_sent_utag_sts_top;
  reg             hd0_cpl_valid_top;
  reg    [0:9]    hd0_cpl_utag_top;
  reg    [0:2]    hd0_cpl_type_top;
  reg    [0:9]    hd0_cpl_size_top;
  reg    [0:9]    hd0_cpl_laddr_top;
  reg    [0:9]    hd0_cpl_byte_count_top;
  reg    [0:1023] hd0_cpl_data_top;
  reg             hd1_sent_utag_valid_top;
  reg    [0:9]    hd1_sent_utag_top;
  reg    [0:2]    hd1_sent_utag_sts_top;
  reg             hd1_cpl_valid_top;
  reg    [0:9]    hd1_cpl_utag_top;
  reg    [0:2]    hd1_cpl_type_top;
  reg    [0:9]    hd1_cpl_size_top;
  reg    [0:9]    hd1_cpl_laddr_top;
  reg    [0:9]    hd1_cpl_byte_count_top;
  reg    [0:1023] hd1_cpl_data_top;

  // Output
  reg             ah_cvalid_top;
  reg    [0:7]    ah_ctag_top;
  reg             ah_ctagpar_top;
  reg    [0:12]   ah_com_top;
  reg             ah_compar_top;
  reg    [0:2]    ah_cabt_top;
  reg    [0:63]   ah_cea_top;
  reg             ah_ceapar_top;
  reg    [0:15]   ah_cch_top;
  reg    [0:11]   ah_csize_top;
  reg    [0:3]    ah_cpagesize_top;
  wire   [0:1023] ah_brdata_top;
  wire   [0:15]   ah_brpar_top;
  wire            ah_brvalid_top;
  wire   [0:7]    ah_brtag_top;
  reg    [0:3]    ah_brlat_top;
  reg             ah_mmack_top;
  reg    [0:63]   ah_mmdata_top;
  reg             ah_mmdatapar_top;
  reg             ah_jdone_top;
  reg             ah_jcack_top;
  reg    [0:63]   ah_jerror_top;
//  reg             ah_jyield_top;
  reg             ah_tbreq_top;
  reg             ah_paren_top;
  reg             d0h_dvalid_top;
  reg    [0:9]    d0h_req_utag_top;
  reg    [0:8]    d0h_req_itag_top;
  reg    [0:2]    d0h_dtype_top;
  reg    [0:9]    d0h_dsize_top;
  reg    [0:1023] d0h_ddata_top;
  reg    [0:5]    d0h_datomic_op_top;
  reg             d0h_datomic_le_top;
  reg             d1h_dvalid_top;
  reg    [0:9]    d1h_req_utag_top;
  reg    [0:8]    d1h_req_itag_top;
  reg    [0:2]    d1h_dtype_top;
  reg    [0:9]    d1h_dsize_top;
  reg    [0:1023] d1h_ddata_top;
  reg    [0:5]    d1h_datomic_op_top;
  reg             d1h_datomic_le_top;

  // Registers
  reg             ah_jrunning_l;
  reg             ha_brvalid;
  reg             ha_bwvalid_l;
  reg             ha_bwvalid;
  reg    [0:7]    ha_bwtag_l;
  reg             ha_bwtagpar_l;
  reg    [0:7]    ha_bwtag;
  reg             ha_bwtagpar;
  reg    [0:1023] ha_bwdata;
  reg    [0:15]   ha_bwpar;
  reg    [0:5]    ha_bwad;
  reg    [0:7]    ha_brtag;
  reg             ha_brtagpar;
  reg    [0:7]    rtag;
  reg             rtagpar;
  reg    [0:8]    rditag;
  reg             rditagpar;
  reg    [0:7]    response;
  reg    [0:8]    response_ext;
  reg    [0:3]    rpagesize;
  reg    [0:1]    rcachestate;
  reg    [0:12]   rcachepos;
  reg    [0:8]    rcredits;
  reg             ha_rvalid;
  reg    [0:7]    ha_rtag;
  reg             ha_rtagpar;
  reg    [0:8]    ha_rditag;
  reg             ha_rditagpar;
  reg    [0:7]    ha_response;
  reg    [0:7]    ha_response_ext;
  reg    [0:3]    ha_rpagesize;
  reg    [0:1]    ha_rcachestate;
  reg    [0:12]   ha_rcachepos;
  reg    [0:8]    ha_rcredits;
  reg             rvalid;
  reg             rvalid_l;
  reg    [0:7]    rtag_l;
  reg             rtagpar_l;
  reg    [0:8]    rditag_l;
  reg             rditagpar_l;
  reg    [0:7]    response_l;
  reg    [0:7]    response_ext_l;
  reg    [0:3]    rpagesize_l;
  reg    [0:1]    rcachestate_l;
  reg    [0:12]   rcachepos_l;
  reg    [0:8]    rcredits_l;
  reg             rvalid_ll;
  reg    [0:7]    rtag_ll;
  reg             rtagpar_ll;
  reg    [0:8]    rditag_ll;
  reg             rditagpar_ll;
  reg    [0:7]    response_ll;
  reg    [0:7]    response_ext_ll;
  reg    [0:3]    rpagesize_ll;
  reg    [0:1]    rcachestate_ll;
  reg    [0:12]   rcachepos_ll;
  reg    [0:8]    rcredits_ll;
  reg    [0:5]    r_wr_ptr;
  reg    [0:5]    r_rd_ptr;
  reg    [0:7]    rtag_array         [0:63];
  reg             rtagpar_array      [0:63];
  reg    [0:8]    rditag_array       [0:63];
  reg             rditagpar_array    [0:63];
  reg    [0:7]    response_array     [0:63];
  reg    [0:7]    response_ext_array [0:63];
  reg    [0:3]    rpagesize_array    [0:63];
  reg    [0:1]    rcachestate_array  [0:63];
  reg    [0:12]   rcachepos_array    [0:63];
  reg    [0:8]    rcredits_array     [0:63];
  reg    [0:5]    bw_wr_ptr;
  reg    [0:5]    bw_rd_ptr;
  reg    [0:5]    bw_rd_ptr_l;
  reg             bwhalf;
  reg    [0:1023] bwdata;
  reg    [0:15]   bwpar;
  reg    [0:1]    bw_active    [0:255];
  reg    [0:5]    br_wr_ptr;
  reg    [0:5]    br_rd_ptr;
  reg    [0:16]   brvalid_delay;
  reg    [0:7]    bwtag_array  [0:63];
  reg             bwtagpar_array[0:63];
  reg    [0:1023] bwdata_array [0:63];
  reg    [0:15]   bwpar_array  [0:63];
  reg    [0:7]    brtag_array  [0:63];
  reg             brtagpar_array[0:63];
  reg    [0:7]    brtag_delay  [0:16];
  reg             brhalf;
//  reg    [0:1023]  brdata_delay;
  reg    [0:7]    brpar_delay;
  reg             hd0_cpl_valid;
  reg    [0:9]    hd0_cpl_utag;
  reg    [0:2]    hd0_cpl_type;
  reg    [0:9]    hd0_cpl_size;
  reg    [0:9]    hd0_cpl_laddr;
  reg    [0:9]    hd0_cpl_byte_count;
  reg    [0:1023] hd0_cpl_data;
  reg             hd1_sent_utag_valid;
  reg    [0:9]    hd1_sent_utag;
  reg    [0:2]    hd1_sent_utag_sts;
  reg             hd1_cpl_valid;
  reg    [0:9]    hd1_cpl_utag;
  reg    [0:2]    hd1_cpl_type;
  reg    [0:9]    hd1_cpl_size;
  reg    [0:9]    hd1_cpl_laddr;
  reg    [0:9]    hd1_cpl_byte_count;
  reg    [0:1023] hd1_cpl_data;
//  reg    [0:15]   hd0_cpl_dpar;

  // Wires
  wire            ah_cvalid;
  wire   [0:7]    ah_ctag;
  wire            ah_ctagpar;
  wire   [0:12]   ah_com;
  wire            ah_compar;
  wire   [0:2]    ah_cabt;
  wire   [0:63]   ah_cea;
  wire            ah_ceapar;
  wire   [0:15]   ah_cch;
  wire   [0:11]   ah_csize;
  wire   [0:3]    ah_cpagesize;
  wire   [0:7]    ha_croom;
  wire            ha_brvalid_ul;
  wire   [0:5]    ha_brad;
  wire   [0:3]    ah_brlat;
  wire   [0:1023] ah_brdata;
  wire   [0:15]   ah_brpar;
  reg             ha_bwvalid_ul;
  wire            ha_mmval;
  wire            ha_mmcfg;
  wire            ha_mmrnw;
  wire            ha_mmdw;
  wire   [0:23]   ha_mmad;
  wire            ha_mmadpar;
  wire   [0:63]   ha_mmdata;
  wire            ha_mmdatapar;
  wire            ah_mmack;
  wire   [0:63]   ah_mmdata;
  wire            ah_mmdatapar;
  wire            ha_jval;
  wire   [0:7]    ha_jcom;
  wire            ha_jcompar;
  wire   [0:63]   ha_jea;
  wire            ha_jeapar;
  wire            ah_jrunning_top;
  wire            ah_jrunning;
  wire            ah_jdone;
  wire            ah_jcack;
  wire   [0:63]   ah_jerror;
//  wire            ah_jyield;
  wire            ah_tbreq;
  wire            ah_paren;
  wire            rvalid_ul;
  reg    [0:185]  ha_reoa;		// UMA : TODO revisit
  wire            d0h_dvalid;
  wire   [0:9]    d0h_req_utag;
  wire   [0:8]    d0h_req_itag;
  wire   [0:2]    d0h_dtype;
  wire   [0:9]    d0h_dsize;
  wire   [0:1023] d0h_ddata;
  wire   [0:5]    d0h_datomic_op;
  wire            d0h_datomic_le;
  wire            d1h_dvalid;
  wire   [0:9]    d1h_req_utag;
  wire   [0:8]    d1h_req_itag;
  wire   [0:2]    d1h_dtype;
  wire   [0:9]    d1h_dsize;
  wire   [0:1023] d1h_ddata;
  wire   [0:5]    d1h_datomic_op;
  wire            d1h_datomic_le;
//  wire   [0:15]   d0h_dpar;
  wire            hd0_sent_utag_valid;
  wire   [0:9]    hd0_sent_utag;
  wire   [0:2]    hd0_sent_utag_sts;

  // Integers

  integer         i;
  reg [0:63]      simulationTime ;
  reg             simulationError;

  // C code interface registration

  initial begin
    ha_pclock <= 0;
    br_wr_ptr <= 0;
    br_rd_ptr <= 0;
    bw_wr_ptr <= 0;
    bw_rd_ptr <= 0;
    r_wr_ptr <= 0;
    r_rd_ptr <= 0;
    ha_jval_top <= 0;
    ha_brvalid_top <= 0;
    ha_bwvalid_top <= 0;
    ha_rvalid_top <= 0;
    ha_croom_top <= 0;
    ha_brtag_top <= 0;
    ha_brtagpar_top <= 0;
    ha_bwtag_top <= 0;
    ha_bwtagpar_top <= 0;
    ha_bwdata_top <= 0;
    ha_bwpar_top <= 0;
    ha_rtag_top <= 0;
    ha_rtagpar_top <= 0;
    ha_rditag_top <= 0;
    ha_rditagpar_top <= 0;
    ha_response_top <= 0;
    ha_response_ext_top <= 0;
    ha_rpagesize_top <= 0;
    ha_rcredits_top <= 9'h01;
    ha_reoa <= 0;
    ha_mmval_top <= 0;
    ha_mmcfg_top <= 0;
    ha_mmrnw_top <= 0;
    ha_mmdw_top <= 0;
    ha_mmad_top <= 0;
    ha_mmadpar_top <= 0;
    ha_mmdata_top <= 0;
    ha_mmdatapar_top <= 0;
    ha_jval_top <= 0;
    ha_jcom_top <= 0;
    ha_jcompar_top <= 0;
    ha_jea_top <= 0;
    ha_jeapar_top <= 0;
    ha_pclock <= 0;
    hd0_sent_utag_valid_top <= 0;
    hd0_sent_utag_top <= 0;
    hd0_sent_utag_sts_top <= 0;
    hd0_cpl_valid_top <= 0;
    hd0_cpl_utag_top <= 0;
    hd0_cpl_type_top <= 0;
    hd0_cpl_size_top <= 0;
    hd0_cpl_laddr_top <= 0;
    hd0_cpl_byte_count_top <= 0;
    hd0_cpl_data_top <= 0;
    hd1_sent_utag_valid_top <= 0;
    hd1_sent_utag_top <= 0;
    hd1_sent_utag_sts_top <= 0;
    hd1_cpl_valid_top <= 0;
    hd1_cpl_utag_top <= 0;
    hd1_cpl_type_top <= 0;
    hd1_cpl_size_top <= 0;
    hd1_cpl_laddr_top <= 0;
    hd1_cpl_byte_count_top <= 0;
    hd1_cpl_data_top <= 0;
    for(i=0; i<64; i++) begin
      bwtag_array[i] <= 0;
      bwtagpar_array[i] <= 0;
      bwdata_array[i] <= 0;
      bwpar_array[i] <= 0;
      brtag_array[i] <= 0;
      brtagpar_array[i] <= 0;
    end
    for(i=0; i<64; i++) begin
      rtag_array[i] <= 0;
      rtagpar_array[i] <= 0;
      rditag_array[i] <= 0;
      rditagpar_array[i] <= 0;
      response_array[i] <= 0;
      response_ext_array[i] <= 0;
      rpagesize_array[i] <= 0;
      rcachestate_array[i] <= 0;
      rcachepos_array[i] <= 0;
      rcredits_array[i] <= 0;
    end
//  hd0_cpl_dpar	<= 0;
    // $afu_init;
     psl_bfm_init();
     brhalf <= 1'b0;
    // $register_clock(ha_pclock);
/*
    $register_control(ha_jval_top, ha_jcom_top, ha_jcompar_top, ha_jea_top,
                      ha_jeapar_top, ah_jrunning_top, ah_jdone_top,
                      ah_jcack_top, ah_jerror_top, ah_brlat_top, ah_jyield,
                      ah_tbreq_top, ah_paren_top);
    $register_mmio(ha_mmval_top, ha_mmcfg_top, ha_mmrnw_top, ha_mmdw_top,
                   ha_mmad_top, ha_mmadpar_top, ha_mmdata_top, ha_mmdatapar_top,
                   ah_mmack_top, ah_mmdata_top, ah_mmdatapar_top);
    $register_command(ha_croom_top, ah_cvalid_top, ah_ctag_top, ah_ctagpar_top,
                      ah_com_top, ah_compar_top, ah_cabt_top,
                      ah_cea_top, ah_ceapar_top, ah_cch_top, ah_csize_top);
    $register_rd_buffer(ha_brvalid_top, ha_brtag_top, ha_brtagpar_top,
                        ah_brdata_top, ah_brpar_top, ah_brvalid_top,
                        ah_brtag_top, ah_brlat_top);
    $register_wr_buffer(ha_bwvalid_top, ha_bwtag_top, ha_bwtagpar_top,
                        ha_bwdata_top, ha_bwpar_top);
    $register_response(ha_rvalid_top, ha_rtag_top, ha_rtagpar_top,
                       ha_response_top, ha_rcredits_top);
*/
  end

  // Clock generation

  always begin
    #2 ha_pclock = !ha_pclock;
  end


  // Passthrough signals

  assign ha_croom     = ha_croom_top;
  assign ha_mmval     = ha_mmval_top;
  assign ha_mmcfg     = ha_mmcfg_top;
  assign ha_mmrnw     = ha_mmrnw_top;
  assign ha_mmdw      = ha_mmdw_top;
  assign ha_mmad      = ha_mmad_top;
  assign ha_mmadpar   = ha_mmadpar_top;
  assign ha_mmdata    = ha_mmdata_top;
  assign ha_mmdatapar = ha_mmdatapar_top;
  assign ha_jval      = ha_jval_top;
  assign ha_jcom      = ha_jcom_top;
  assign ha_jcompar   = ha_jcompar_top;
  assign ha_jea       = ha_jea_top;
  assign ha_jeapar    = ha_jeapar_top;
  assign hd0_sent_utag_valid    = hd0_sent_utag_valid_top;
  assign hd0_sent_utag    	= hd0_sent_utag_top;
  assign hd0_sent_utag_sts    	= hd0_sent_utag_sts_top;
  assign hd0_cpl_valid    	= hd0_cpl_valid_top;
  assign hd0_cpl_utag    	= hd0_cpl_utag_top;
  assign hd0_cpl_type    	= hd0_cpl_type_top;
  assign hd0_cpl_size    	= hd0_cpl_size_top;
  assign hd0_cpl_laddr    	= hd0_cpl_laddr_top;
  assign hd0_cpl_byte_count    	= hd0_cpl_byte_count_top;
  assign hd0_cpl_data    	= hd0_cpl_data_top;
  assign hd1_sent_utag_valid    = hd1_sent_utag_valid_top;
  assign hd1_sent_utag    	= hd1_sent_utag_top;
  assign hd1_sent_utag_sts    	= hd1_sent_utag_sts_top;
  assign hd1_cpl_valid    	= hd1_cpl_valid_top;
  assign hd1_cpl_utag    	= hd1_cpl_utag_top;
  assign hd1_cpl_type    	= hd1_cpl_type_top;
  assign hd1_cpl_size    	= hd1_cpl_size_top;
  assign hd1_cpl_laddr    	= hd1_cpl_laddr_top;
  assign hd1_cpl_byte_count    	= hd1_cpl_byte_count_top;
  assign hd1_cpl_data    	= hd1_cpl_data_top;

  always @ ( ha_pclock ) begin
    simulationTime = $time;
    set_simulation_time(simulationTime);
//    $display("%d : Calling to C ", simulationTime);
    psl_bfm( ha_pclock, 
             ha_jval_top, 
             ha_jcom_top, 
             ha_jcompar_top, 
             ha_jea_top,
	     ha_jeapar_top, 
             ah_jrunning_top,  
             ah_jdone_top,
	     ah_jcack_top, 
             ah_jerror_top, 
             ah_brlat_top,  
//             ah_jyield,
	     ah_tbreq_top, 
             ah_paren_top, 
             ha_mmval_top,
             ha_mmcfg_top, 
             ha_mmrnw_top, 
             ha_mmdw_top,
             ha_mmad_top, 
             ha_mmadpar_top, 
             ha_mmdata_top, 
             ha_mmdatapar_top,
             ah_mmack_top, 
             ah_mmdata_top, 
             ah_mmdatapar_top,
             ha_croom_top,
             ah_cvalid_top, 
             ah_ctag_top, 
             ah_ctagpar_top, 
             ah_com_top, 
             ah_compar_top, 
             ah_cabt_top, 
             ah_cea_top, 
             ah_ceapar_top, 
             ah_cch_top, 
             ah_csize_top, 
             ah_cpagesize_top, 
             ha_brvalid_top, 
             ha_brtag_top, 
             ha_brtagpar_top, 
             ah_brdata_top, 
             ah_brpar_top, 
             ah_brvalid_top, 
             ah_brtag_top,
             ha_bwvalid_top, 
             ha_bwtag_top, 		// 8 bits
             ha_bwtagpar_top,
             ha_bwdata_top, 		// 1024 bits
             ha_bwpar_top,	// 16 bits
             ha_rvalid_top, 
             ha_rtag_top, 		// 8 bits
             ha_rtagpar_top,
             ha_rditag_top,		// 9 bits
             ha_rditagpar_top,
             ha_response_top, 		// 8 bits
             ha_response_ext_top, 	// 8 bits
             ha_rpagesize_top,	 	// 4 bits
             ha_rcachestate_top, 	// 2 bits
             ha_rcachepos_top, 		// 13 bits
             ha_rcredits_top,		// 9 bits
             d0h_dvalid_top, 		// DMA Port 0
             d0h_req_utag_top, 
             d0h_req_itag_top, 
             d0h_dtype_top, 
             d0h_dsize_top, 
             d0h_ddata_top, 
             d0h_datomic_op_top, 
             d0h_datomic_le_top, 
	     hd0_sent_utag_valid_top, 
	     hd0_sent_utag_top, 
	     hd0_sent_utag_sts_top, 
	     hd0_cpl_valid_top,  
	     hd0_cpl_utag_top,  
	     hd0_cpl_type_top,  
	     hd0_cpl_size_top,  
	     hd0_cpl_laddr_top,  
	     hd0_cpl_byte_count_top,  
	     hd0_cpl_data_top,  
             d1h_dvalid_top, 		// DMA Port 1
             d1h_req_utag_top, 
             d1h_req_itag_top, 
             d1h_dtype_top, 
             d1h_dsize_top, 
             d1h_ddata_top, 
             d1h_datomic_op_top, 
             d1h_datomic_le_top, 
	     hd1_sent_utag_valid_top, 
	     hd1_sent_utag_top, 
	     hd1_sent_utag_sts_top, 
	     hd1_cpl_valid_top,  
	     hd1_cpl_utag_top,  
	     hd1_cpl_type_top,  
	     hd1_cpl_size_top,  
	     hd1_cpl_laddr_top,  
	     hd1_cpl_byte_count_top,  
	     hd1_cpl_data_top
             );
  end

  always @ (negedge ha_pclock) begin
    get_simuation_error(simulationError);
  end

  always @ (posedge ha_pclock) begin
    ah_jrunning_l <= ah_jrunning;
    if(simulationError)
      $finish;
//      $stop;
  end

  assign ah_jrunning_top = ah_jrunning_l;

  // Latch top level signals

  always @ (posedge ha_pclock) begin
    ah_ctag_top <= ah_ctag;
    ah_ctagpar_top <= ah_ctagpar;
    ah_com_top <= ah_com;
    ah_compar_top <= ah_compar;
    ah_cabt_top <= ah_cabt;
    ah_cea_top <= ah_cea;
    ah_ceapar_top <= ah_ceapar;
    ah_cch_top <= ah_cch;
    ah_csize_top <= ah_csize;
    ah_cpagesize_top <= ah_cpagesize;
    ah_mmdata_top <= ah_mmdata;
    ah_mmdatapar_top <= ah_mmdatapar;
    ah_jerror_top <= ah_jerror;
    ah_jdone_top <= ah_jdone;
    ah_brlat_top <= ah_brlat;
//    ah_jyield_top <= ah_jyield;
    ah_tbreq_top <= ah_tbreq;
    ah_paren_top <= ah_paren;
    ah_cvalid_top <= ah_cvalid;
    ah_mmack_top <= ah_mmack;
    ah_jcack_top <= ah_jcack;
    d0h_dvalid_top <= d0h_dvalid;
    d0h_req_utag_top <= d0h_req_utag;
    d0h_req_itag_top <= d0h_req_itag;
    d0h_dtype_top <= d0h_dtype;
    d0h_dsize_top <= d0h_dsize;
    d0h_ddata_top <= d0h_ddata;
    d0h_datomic_op_top <= d0h_datomic_op;
    d0h_datomic_le_top <= d0h_datomic_le;
    d1h_dvalid_top <= d1h_dvalid;
    d1h_req_utag_top <= d1h_req_utag;
    d1h_req_itag_top <= d1h_req_itag;
    d1h_dtype_top <= d1h_dtype;
    d1h_dsize_top <= d1h_dsize;
    d1h_ddata_top <= d1h_ddata;
    d1h_datomic_op_top <= d1h_datomic_op;
    d1h_datomic_le_top <= d1h_datomic_le;
  end

  // Breakpoint output, need at least 1 output or Quartus will optimize away
  // and fail to compile.

  assign breakpoint = ah_mmack_top | ah_cvalid_top | ah_brvalid_top |
                      ah_jdone | ah_jcack | (ah_jrunning & !ah_jrunning_l);

  // Buffer write

  always @ (posedge ha_pclock) begin
    for (i = 0; i < 256; i = i + 1) begin
      if (ha_bwvalid_top & (i==ha_bwtag_top))
        bw_active[i] <= bw_active[i] + 1;
       else if (bwhalf & (i==ha_bwtag_l))
         bw_active[i] <= bw_active[i] - 1;
      else if (bw_wr_ptr == bw_rd_ptr)
        bw_active[i] <= 1'b0;
      else
        bw_active[i] <= bw_active[i];
    end
  end

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_top)
      bw_wr_ptr <= bw_wr_ptr+6'h01;
    else
      bw_wr_ptr <= bw_wr_ptr;
  end

  always @ (posedge ha_pclock) begin
     if (ha_bwvalid_l & !bwhalf)
       bw_rd_ptr <= bw_rd_ptr+6'h01;
     else
      bw_rd_ptr <= bw_rd_ptr;
  end

  always @ (posedge ha_pclock)
    bw_rd_ptr_l <= bw_rd_ptr;

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_top)
      bwtag_array[bw_wr_ptr] <= ha_bwtag_top;
  end

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_top)
      bwtagpar_array[bw_wr_ptr] <= ha_bwtagpar_top;
  end

  always @ (posedge ha_pclock)
    ha_bwvalid_ul <= ha_bwvalid_top;

//  assign ha_bwvalid_ul = (bw_rd_ptr==bw_wr_ptr) ? 1'b0 : 1'b1;

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_ul)
      ha_bwtag_l <= bwtag_array[bw_rd_ptr];
    else
      ha_bwtag_l <= 8'b0;
  end

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_ul)
      ha_bwtagpar_l <= bwtagpar_array[bw_rd_ptr];
    else
      ha_bwtagpar_l <= 1'b1;
  end

  always @ (posedge ha_pclock)
    ha_bwtag <= ha_bwtag_l;

  always @ (posedge ha_pclock)
    ha_bwtagpar <= ha_bwtagpar_l;

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_top)
      bwdata_array[bw_wr_ptr] <= ha_bwdata_top;
  end

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_ul)
      bwdata <= bwdata_array[bw_rd_ptr];
  end

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_top)
      bwpar_array[bw_wr_ptr] <= ha_bwpar_top;
  end

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_ul)
      // bwpar <= bwpar_array[bw_rd_ptr_l];  // this is the p8 method because parity lags data by one cycle
      bwpar <= bwpar_array[bw_rd_ptr];  // this the p9 method because parity and data are coincident
  end

  always @ (posedge ha_pclock)
    ha_bwvalid_l <= ha_bwvalid_ul;

  always @ (posedge ha_pclock)
    ha_bwvalid <= ha_bwvalid_l;

  always @ (posedge ha_pclock) begin
    if (ha_bwvalid_l & !bwhalf)
      bwhalf <= 1;
    else
      bwhalf <= 0;
  end

  always @ (posedge ha_pclock)
//    ha_bwad <= {5'b0, bwhalf};
    ha_bwad <= {6'b0};

  always @ (posedge ha_pclock) begin
    if (!bwhalf)
      ha_bwdata <= bwdata[0:1023];
    else
      ha_bwdata <= bwdata[0:1023];
  end

  always @ (posedge ha_pclock) begin
    if (bwhalf)
      ha_bwpar <= bwpar[0:15];
    else
     ha_bwpar <= bwpar[0:15];
  end

  // Buffer read

  always @ (posedge ha_pclock) begin
    if (ha_brvalid_top)
      br_wr_ptr <= br_wr_ptr+6'h01;
    else
      br_wr_ptr <= br_wr_ptr;
  end

  always @ (posedge ha_pclock) begin
    if (ha_brvalid & !brhalf)
      br_rd_ptr <= br_rd_ptr+6'h01;
    else
      br_rd_ptr <= br_rd_ptr;
  end

  always @ (posedge ha_pclock) begin
    for (i = 0; i <= 16; i = i + 1) begin
      if (i == ah_brlat+1) begin
        brvalid_delay[i] <= ha_brvalid  & !brhalf;
        brtag_delay[i] <= ha_brtag;
      end else if (i == 16) begin
        brvalid_delay[16] <= 1'b0;
        brtag_delay[16] <= 8'h00;
      end else begin
        brvalid_delay[i] <= brvalid_delay[i+1];
        brtag_delay[i] <= brtag_delay[i+1];
      end
    end
  end

  always @ (posedge ha_pclock) begin
    if (ha_brvalid_top)
      brtag_array[br_wr_ptr] <= ha_brtag_top;
  end

  always @ (posedge ha_pclock) begin
    if (ha_brvalid_top)
      brtagpar_array[br_wr_ptr] <= ha_brtagpar_top;
  end

  assign ha_brvalid_ul = (br_rd_ptr==br_wr_ptr) ? 1'b0 : 1'b1;

  always @ (posedge ha_pclock) begin
    if (ha_brvalid_ul)
      ha_brtag <= brtag_array[br_rd_ptr];
  end

  always @ (posedge ha_pclock) begin
    if (ha_brvalid_ul)
      ha_brtagpar <= brtagpar_array[br_rd_ptr];
  end

  always @ (posedge ha_pclock) begin
    if (br_rd_ptr==br_wr_ptr)
      ha_brvalid <= 1'b0;
    else
      ha_brvalid <= 1'b1;
  end
/*
  always @ (posedge ha_pclock) begin
    if (ha_brvalid & !brhalf)
      brhalf <= 1'b1;
    else
      brhalf <= 1'b0;
  end
*/
//  assign ha_brad = {5'b0, brhalf};
  assign ha_brad = {6'b0};
 
  always @ (posedge ha_pclock) begin
//    brdata_delay <= ah_brdata;
  end

  always @ (posedge ha_pclock) begin
    brpar_delay <= ah_brpar;
  end

//  assign ah_brdata_top = {brdata_delay, ah_brdata};
  assign ah_brdata_top = ah_brdata;
//  assign ah_brpar_top = {brpar_delay, ah_brpar};
  assign ah_brpar_top =  ah_brpar;
  assign ah_brvalid_top = brvalid_delay[0];
  assign ah_brtag_top = brtag_delay[0];

  // Response delay

  always @ (posedge ha_pclock) begin
    if (ha_rvalid_top)
      r_wr_ptr <= r_wr_ptr+6'h01;
    else
      r_wr_ptr <= r_wr_ptr;
  end

  assign rvalid_ul = (r_wr_ptr!=r_rd_ptr) &
                     (bw_active[rtag_array[r_rd_ptr]]==0);

  always @ (posedge ha_pclock) begin
    if (rvalid_ul)
      r_rd_ptr <= r_rd_ptr+6'h01;
    else
      r_rd_ptr <= r_rd_ptr;
  end

  always @ (posedge ha_pclock) begin
    if (ha_rvalid_top) begin
      rtag_array[r_wr_ptr] 		<= ha_rtag_top;
      rtagpar_array[r_wr_ptr] 		<= ha_rtagpar_top;
      rditag_array[r_wr_ptr] 		<= ha_rditag_top;
      rditagpar_array[r_wr_ptr]		<= ha_rditagpar_top;
      response_array[r_wr_ptr] 		<= ha_response_top;
      response_ext_array[r_wr_ptr] 	<= ha_response_ext_top;
      rpagesize_array[r_wr_ptr]	 	<= ha_rpagesize_top;
      rcachestate_array[r_wr_ptr] 	<= ha_rcachestate_top;
      rcachepos_array[r_wr_ptr] 	<= ha_rcachepos_top;
      rcredits_array[r_wr_ptr] 		<= ha_rcredits_top;
    end
  end

  always @ (posedge ha_pclock) begin
    if (rvalid_ul) begin
      rtag 		<= rtag_array[r_rd_ptr];
      rtagpar 		<= rtagpar_array[r_rd_ptr];
      rditag 		<= rditag_array[r_rd_ptr];
      rditagpar 	<= rditagpar_array[r_rd_ptr];
      response 		<= response_array[r_rd_ptr];
      response_ext 	<= response_ext_array[r_rd_ptr];
      rpagesize 	<= rpagesize_array[r_rd_ptr];
      rcachestate 	<= rcachestate_array[r_rd_ptr];
      rcachepos 	<= rcachepos_array[r_rd_ptr];
      rcredits 		<= rcredits_array[r_rd_ptr];
    end
  end

  always @ (posedge ha_pclock) begin
    rvalid <= rvalid_ul;
    rvalid_l <= rvalid;
    rtag_l <= rtag;
    rtagpar_l <= rtagpar;
    rditag_l <= rditag;
    rditagpar_l <= rditagpar;
    response_l <= response;
    response_ext_l <= response_ext;
    rpagesize_l <= rpagesize;
    rcachestate_l <= rcachestate;
    rcachepos_l <= rcachepos;
    rcredits_l <= rcredits;
    rvalid_ll <= rvalid_l;
    rtag_ll <= rtag_l;
    rtagpar_ll <= rtagpar_l;
    rditag_ll <= rditag_l;
    rditagpar_ll <= rditagpar_l;
    response_ll <= response_l;
    response_ext_ll <= response_ext_l;
    rpagesize_ll <= rpagesize_l;
    rcachestate_ll <= rcachestate_l;
    rcachepos_ll <= rcachepos_l;
    rcredits_ll <= rcredits_l;
    ha_rvalid <= rvalid_ll;
    ha_rtag <= rtag_ll;
    ha_rtagpar <= rtagpar_ll;
    ha_rditag <= rditag_ll;
    ha_rditagpar <= rditagpar_ll;
    ha_response <= response_ll;
    ha_response_ext <= response_ext_ll;
    ha_rpagesize <= rpagesize_ll;
//    ha_rcachestate <= rcachestate_ll;
    ha_rcachestate <= 0;			// Since this is a reserved signal, driving it to '0' as of now	:TODO: UMA will update, if there is a definition
//    ha_rcachepos <= rcachepos_ll;
    ha_rcachepos <= 0;			// Since this is a reserved signal, driving it to '0' as of now	:TODO: UMA will update, if there is a definition
//    ha_rcredits <= rcredits_ll;
    ha_rcredits <= 9'h1;		// Defined as reserved, but requires a static value of 9'b000000001 to indicate 1 credit is always
  end

  // AFU instance

  mcp_top a0 (
    // Command interface
    .ah_cvalid(ah_cvalid),
    .ah_ctag(ah_ctag),
    .ah_ctagpar(ah_ctagpar),
    .ah_com(ah_com),
    .ah_compar(ah_compar),
    .ah_cabt(ah_cabt),
    .ah_cea(ah_cea),
    .ah_ceapar(ah_ceapar),
    .ah_cch(ah_cch),
    .ah_csize(ah_csize),
    .ah_cpagesize(ah_cpagesize),
    .ha_croom(ha_croom),
    // Buffer interface
    .ha_brvalid(ha_brvalid),
    .ha_brtag(ha_brtag),
    .ha_brtagpar(ha_brtagpar),
    .ha_brad(ha_brad),				// UMA - TODO - should revisit
    .ah_brlat(ah_brlat),
    .ah_brdata(ah_brdata),
    .ah_brpar(ah_brpar),
    .ha_bwvalid(ha_bwvalid),
    .ha_bwtag(ha_bwtag),
    .ha_bwtagpar(ha_bwtagpar),
    .ha_bwad(ha_bwad),
    .ha_bwdata(ha_bwdata),
    .ha_bwpar(ha_bwpar),
    // Response interface
    .ha_rvalid(ha_rvalid),
    .ha_rtag(ha_rtag),
    .ha_rtagpar(ha_rtagpar),
    .ha_rditag(ha_rditag),
    .ha_rditagpar(ha_rditagpar),
    .ha_response(ha_response),
    .ha_response_ext(ha_response_ext),
    .ha_rpagesize(ha_rpagesize),
    .ha_rcredits(ha_rcredits),
    .ha_rcachestate(ha_rcachestate),
    .ha_rcachepos(ha_rcachepos),
//    .ha_reoa(ha_reoa),	- mcp004 does not seem to have this port
    // MMIO interface
    .ha_mmval(ha_mmval),
    .ha_mmcfg(ha_mmcfg),
    .ha_mmrnw(ha_mmrnw),
    .ha_mmdw(ha_mmdw),
    .ha_mmad(ha_mmad),
    .ha_mmadpar(ha_mmadpar),
    .ha_mmdata(ha_mmdata),
    .ha_mmdatapar(ha_mmdatapar),
    .ah_mmack(ah_mmack),
    .ah_mmdata(ah_mmdata),
    .ah_mmdatapar(ah_mmdatapar),
    // Control interface
    .ha_jval(ha_jval),
    .ha_jcom(ha_jcom),
    .ha_jcompar(ha_jcompar),
    .ha_jea(ha_jea),
    .ha_jeapar(ha_jeapar),
    .ah_jrunning(ah_jrunning),
    .ah_jdone(ah_jdone),
    .ah_jcack(ah_jcack),
    .ah_jerror(ah_jerror),
//    .ah_jyield(ah_jyield),	- mcp004 does not seem to have this port
    .ah_tbreq(ah_tbreq),
    .ah_paren(ah_paren),
    .ha_pclock(ha_pclock),
    // DMA 0 Req interface
    .d0h_dvalid(d0h_dvalid),
    .d0h_req_utag(d0h_req_utag),
    .d0h_req_itag(d0h_req_itag),
    .d0h_dtype(d0h_dtype),
    .d0h_dsize(d0h_dsize),
    .d0h_ddata(d0h_ddata),
    .d0h_datomic_op(d0h_datomic_op),				
    .d0h_datomic_le(d0h_datomic_le),		
//    .d0h_dpar(d0h_dpar),
    // DMA 0 Sent interface
    .hd0_sent_utag_valid(hd0_sent_utag_valid),
    .hd0_sent_utag(hd0_sent_utag),
    .hd0_sent_utag_sts(hd0_sent_utag_sts),
    // DMA 0 CPL interface
    .hd0_cpl_valid(hd0_cpl_valid),
    .hd0_cpl_utag(hd0_cpl_utag),
    .hd0_cpl_type(hd0_cpl_type),
    .hd0_cpl_size(hd0_cpl_size),
    .hd0_cpl_laddr(hd0_cpl_laddr),
    .hd0_cpl_byte_count(hd0_cpl_byte_count),
    .hd0_cpl_data(hd0_cpl_data),
//    .hd0_cpl_dpar(hd0_cpl_dpar)
    // DMA 1 Req interface
    .d1h_dvalid(d1h_dvalid),
    .d1h_req_utag(d1h_req_utag),
    .d1h_req_itag(d1h_req_itag),
    .d1h_dtype(d1h_dtype),
    .d1h_dsize(d1h_dsize),
    .d1h_ddata(d1h_ddata),
    .d1h_datomic_op(d1h_datomic_op),				
    .d1h_datomic_le(d1h_datomic_le),			
    // DMA 1 Sent interface
    .hd1_sent_utag_valid(hd1_sent_utag_valid),
    .hd1_sent_utag(hd1_sent_utag),
    .hd1_sent_utag_sts(hd1_sent_utag_sts),
    // DMA 1 CPL interface
    .hd1_cpl_valid(hd1_cpl_valid),
    .hd1_cpl_utag(hd1_cpl_utag),
    .hd1_cpl_type(hd1_cpl_type),
    .hd1_cpl_size(hd1_cpl_size),
    .hd1_cpl_laddr(hd1_cpl_laddr),
    .hd1_cpl_byte_count(hd1_cpl_byte_count),
    .hd1_cpl_data(hd1_cpl_data)
  );

endmodule
